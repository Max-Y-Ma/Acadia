// Configuration for UVM Testbench for RISCV Pipeline CPU
`define NUM_TEST (500000)
`define NOP_INSTR (32'h13)