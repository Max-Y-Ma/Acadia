adsfasd
  adsf