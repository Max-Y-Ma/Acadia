module core (

);


endmodule : core