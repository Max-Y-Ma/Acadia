// Toggle Test Types
// `define CONSTRAINED_RANDOM  // Comment out for directed tests

`ifdef CONSTRAINED_RANDOM
    `include "cpu_pkg.svh"
`endif

module top_tb;
    timeunit 1ps;
    timeprecision 1ps;

    // UVM Imports
    `ifdef CONSTRAINED_RANDOM
        import uvm_pkg::*;
        `include "uvm_macros.svh"
    `endif

    // Clock Generation
    `define CLK_HALF_PERIOD (5)
    bit clk;
    always #(`CLK_HALF_PERIOD) clk = ~clk;

    bit rst;

    // Memory Interface
    mem_itf mem_itf_i(.clk(clk), .rst(rst));
    mem_itf mem_itf_d(.clk(clk), .rst(rst));

    // Monitor Interface
    mon_itf mon_itf(.*);    
    monitor monitor(.itf(mon_itf));

    // Test Suite
    `ifdef CONSTRAINED_RANDOM
        initial begin
            // UVM Constrained Random Tests
            uvm_config_db #(virtual mem_itf)::set(null, "*", "mem_itf_i", mem_itf_i);
            uvm_config_db #(virtual mem_itf)::set(null, "*", "mem_itf_d", mem_itf_d);
            run_test();
        end
    `else
        // Memory Types for Directed Test
        // magic_dual_port mem(.itf_i(mem_itf_i), .itf_d(mem_itf_d));
        ordinary_dual_port mem(.itf_i(mem_itf_i), .itf_d(mem_itf_d));
    `endif

    // DUT Instantiation
    cpu dut(
        .clk            (clk),
        .rst            (rst),

        // Instruction Memory Port
        .imem_addr      (mem_itf_i.addr),
        .imem_rmask     (mem_itf_i.rmask),
        .imem_rdata     (mem_itf_i.rdata),
        .imem_resp      (mem_itf_i.resp),

        // Data Memory Port
        .dmem_addr      (mem_itf_d.addr),
        .dmem_rmask     (mem_itf_d.rmask),
        .dmem_wmask     (mem_itf_d.wmask),
        .dmem_rdata     (mem_itf_d.rdata),
        .dmem_wdata     (mem_itf_d.wdata),
        .dmem_resp      (mem_itf_d.resp)
    );

    // Monitor Interface DUT Wiring
    `include "../../hvl/rvfi_reference.svh"

    // Waveform Dumpfiles and Reset
    initial begin
        $fsdbDumpfile("dump.fsdb");
        $fsdbDumpvars(0, "+all");
        rst = 1'b1;
        repeat (2) @(posedge clk);
        rst <= 1'b0;
    end

    // End Condition
    int timeout_cycles = 10000000;
    always @(posedge clk) begin
        if (mon_itf.halt) begin
            $finish;
        end
        if (timeout_cycles == 0) begin
            $error("TB Error: Timed out");
            $finish;
        end
        if (mon_itf.error != 0) begin
            repeat (5) @(posedge clk);
            $finish;
        end
        if (mem_itf_i.error != 0) begin
            repeat (5) @(posedge clk);
            $finish;
        end
        if (mem_itf_d.error != 0) begin
            repeat (5) @(posedge clk);
            $finish;
        end
        timeout_cycles <= timeout_cycles - 1;
    end
endmodule : top_tb
